module and_gate (a, b, o);

input a;
input b;
output o;

assign o = a & b;

endmodule